module pipe_MIPS32 (clk1,clk2);
     input clk1,clk2;//two-phase clock
//defining sub-stage variables at different stages
reg [31:0] PC,IF_ID_IR,IF_ID_NPC;
reg [31:0] ID_EX_IR,ID_EX_NPC,ID_EX_A,ID_EX_B,ID_EX_Imm;
reg [2:0] ID_EX_type,EX_MEM_type,MEM_WB_type;
reg [31:0] EX_MEM_IR,EX_MEM_ALUout,EX_MEM_B
reg        EX_MEM_cond;
reg [31:0] MEM_WB_IR,MEM_WB_ALUout,MEM_WB_LMD;

reg [31:0] Reg [0:31];//register bank (32x32)
reg [31:0] Mem [0:1023];//1025x32 memory

parameter ADD=6'b000000, SUB=6'b000001, AND=6'b000010, OR=6'b000011, SLT=6'b000100, MUL=6'b000101,HLT=6'b111111,LW=6'b001000,SW=6'b001001,ADDI=6'b001010,SUBI=6'b001011,SLTI=6'b001100,BNEQZ=6'b001101,BEQZ=6'b001110;
parameter RR_ALU=3'b000, RM_ALU=3'b001, LOAD=3'b010, STORE=3'b011, BRANCH=3'b100, HALT=3'b101;


reg HALTED;
     //Set after HLT instruction is completed(in WB stage)
reg TAKEN_BRANCH;
     //Required to disable instructions after branch

//IF Stage
always @(posedge clk1)                                  // IF Stage
if (HALTED == 0)
begin
  if (((EX_MEM_IR[31:26] == BEQZ) && (EX_MEM_cond == 1)) || ((EX_MEM_IR[31:26] == BNEQZ) && (EX_MEM_cond == 0)))
     begin
          IF_ID_IR      <= #2 Mem[EX_MEM_ALUout];
          TAKEN_BRANCH  <= #2 1'b1;
          IF_ID_NPC     <= #2 EX_MEM_ALUout + 1;
          PC            <= #2 EX_MEM_ALUout + 1;
     end
  else
     begin
          IF_ID_IR      <= #2 Mem[PC];
          IF_ID_NPC     <= #2 PC + 1;
          PC            <= #2 PC + 1;
     end
end





endmodule